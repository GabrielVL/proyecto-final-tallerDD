`timescale 1ns/1ps

module ram_tb;
    logic [14:0] address_a, address_b;
    logic clock;
    logic [7:0] data_a, data_b;
    logic wren_a, wren_b;
    logic [7:0] q_a, q_b;

    ram ram_inst (
        .address_a(address_a),
        .address_b(address_b),
        .clock(clock),
        .data_a(data_a),
        .data_b(data_b),
        .wren_a(wren_a),
        .wren_b(wren_b),
        .q_a(q_a),
        .q_b(q_b)
    );

    initial begin
        clock = 0;
        forever #5 clock = ~clock;
    end

    initial begin
        address_a = 0;
        address_b = 0;
        data_a = 0;
        data_b = 0;
        wren_a = 0;
        wren_b = 0;
        #20;
        $display("Time=%t q_a=%h q_b=%h", $time, q_a, q_b);
        $finish;
    end
endmodule